full_adder_inst : full_adder PORT MAP (
		cin	 => cin_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		cout	 => cout_sig,
		result	 => result_sig
	);
