library verilog;
use verilog.vl_types.all;
entity UART_RX_vlg_vec_tst is
end UART_RX_vlg_vec_tst;
