-------------------------------------------------------------------------------
-- Project     : Audio_Synth
-- Description : Constants and LUT for audio filters
--
--
-------------------------------------------------------------------------------
--
-- Change History
-- Date     |Name      |Modification
------------|----------|-------------------------------------------------------
-- 26.03.18 | dqtm     | file created for EA-999 demo
-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
-- Package  Declaration
-------------------------------------------------------------------------------
-- Include in Design of filter blocks, using  :
--   use work.audio_filter_pkg.all;
-------------------------------------------------------------------------------
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

package audio_filter_pkg is

    --constant N_CUM:					natural :=19; 			-- number of bits in phase cumulator phicum_reg
	--constant N_AUDIO :				natural := 16;			-- Audio Paralell Bus width

    -------------------------------------------------------------------------------
	-- CONSTANT & TYPES FOR FIR 
	-------------------------------------------------------------------------------
    constant N_RESOL_TAP:			natural := 32;  		-- resolution of each position on tap-line (storing MAC outputs)
    constant N_LUT:					natural := 255;  		-- length of LUT = 255
	constant N_addr_LUT:			natural := 8; 			-- number of bits to address LUT (for index)
	
    constant N_RESOL_COEFF:			natural := 16;			-- Attention: 1 bit reserved for sign, FIR-coeffs use 12-bits
															-- range : [-2^15; +(2^15)-1] = [-32768 ; +32767]
															-- but from Matlab file expect scaling fitting in the
															-- range : [-2^11; +(2^11)-1] = [-2048 ; +2047]
    subtype  t_fir_range is integer range -(2**(N_RESOL_COEFF-1)) to (2**(N_RESOL_COEFF-1))-1;
	type     t_lut_fir is array (0 to N_LUT-1) of t_fir_range;


	constant LUT_FIR_LPF_200Hz : t_lut_fir :=(
	-14,-15,-19,-25,-34,-45,-58,-73,-90,-109,-129,-149,-170,-189,-208,
	-226,-241,-253,-263,-269,-272,-273,-273,-273,-272,-270,-268,-265,-262,
	-257,-252,-247,-240,-233,-225,-216,-207,-197,-186,-174,-161,-147,-133,
	-118,-102,-85,-67,-49,-29,-9,12,33,56,79,103,128,154,180,207,235,264,
	293,322,353,384,415,447,480,513,547,580,615,649,685,720,755,791,827,
	863,900,936,972,1009,1045,1081,1118,1154,1189,1225,1260,1295,1330,
	1364,1398,1431,1464,1496,1528,1559,1589,1619,1648,1676,1703,1730,1755,
	1780,1804,1827,1848,1869,1889,1908,1925,1942,1957,1971,1984,1996,2007,
	2016,2024,2031,2037,2041,2044,2046,2047,2046,2044,2041,2037,2031,2024,
	2016,2007,1996,1984,1971,1957,1942,1925,1908,1889,1869,1848,1827,1804,
	1780,1755,1730,1703,1676,1648,1619,1589,1559,1528,1496,1464,1431,1398,
	1364,1330,1295,1260,1225,1189,1154,1118,1081,1045,1009,972,936,900,
	863,827,791,755,720,685,649,615,580,547,513,480,447,415,384,353,322,
	293,264,235,207,180,154,128,103,79,56,33,12,-9,-29,-49,-67,-85,-102,
	-118,-133,-147,-161,-174,-186,-197,-207,-216,-225,-233,-240,-247,-252,
	-257,-262,-265,-268,-270,-272,-273,-273,-273,-272,-269,-263,-253,-241,
	-226,-208,-189,-170,-149,-129,-109,-90,-73,-58,-45,-34,-25,-19,-15,-14
	);
	
	constant LUT_FIR_LPF_400Hz : t_lut_fir :=(
	8,9,11,15,21,27,35,45,55,66,77,89,99,109,118,124,129,132,132,130,125,
	119,112,104,95,86,75,64,52,40,26,12,-2,-17,-33,-49,-65,-82,-99,-116,
	-134,-151,-168,-185,-202,-219,-235,-251,-266,-281,-295,-308,-320,-330,
	-340,-349,-356,-362,-366,-369,-370,-370,-367,-363,-357,-349,-339,-327,
	-312,-296,-278,-257,-234,-209,-182,-153,-121,-88,-52,-15,25,66,110,
	155,201,250,300,351,404,458,513,569,625,683,741,799,858,917,976,1034,
	1093,1151,1208,1264,1320,1374,1428,1480,1530,1579,1626,1671,1714,1755,
	1793,1830,1863,1894,1923,1948,1971,1991,2008,2022,2033,2041,2045,2047,
	2045,2041,2033,2022,2008,1991,1971,1948,1923,1894,1863,1830,1793,1755,
	1714,1671,1626,1579,1530,1480,1428,1374,1320,1264,1208,1151,1093,1034,
	976,917,858,799,741,683,625,569,513,458,404,351,300,250,201,155,110,
	66,25,-15,-52,-88,-121,-153,-182,-209,-234,-257,-278,-296,-312,-327,
	-339,-349,-357,-363,-367,-370,-370,-369,-366,-362,-356,-349,-340,-330,
	-320,-308,-295,-281,-266,-251,-235,-219,-202,-185,-168,-151,-134,-116,
	-99,-82,-65,-49,-33,-17,-2,12,26,40,52,64,75,86,95,104,112,119,125,
	130,132,132,129,124,118,109,99,89,77,66,55,45,35,27,21,15,11,9,8
	);

	constant LUT_FIR_LPF_800Hz : t_lut_fir :=(
	4,4,6,8,11,15,20,25,30,36,40,44,47,48,48,45,40,33,25,15,3,-8,-20,
	-32,-45,-57,-69,-80,-90,-100,-109,-116,-122,-126,-129,-130,-129,
	-126,-121,-115,-106,-96,-83,-69,-54,-37,-19,0,20,41,61,82,102,122,
	140,158,174,188,199,209,216,220,220,218,213,204,192,177,158,136,
	111,84,54,22,-12,-47,-84,-121,-158,-194,-230,-264,-296,-326,-352,
	-375,-394,-408,-416,-420,-417,-408,-393,-371,-342,-306,-263,-213,
	-157,-94,-24,52,133,219,310,405,504,605,708,813,918,1023,1126,1228,
	1327,1422,1513,1599,1679,1753,1819,1878,1929,1971,2004,2028,2042,
	2047,2042,2028,2004,1971,1929,1878,1819,1753,1679,1599,1513,1422,
	1327,1228,1126,1023,918,813,708,605,504,405,310,219,133,52,-24,-94,
	-157,-213,-263,-306,-342,-371,-393,-408,-417,-420,-416,-408,-394,
	-375,-352,-326,-296,-264,-230,-194,-158,-121,-84,-47,-12,22,54,84,
	111,136,158,177,192,204,213,218,220,220,216,209,199,188,174,158,
	140,122,102,82,61,41,20,0,-19,-37,-54,-69,-83,-96,-106,-115,-121,
	-126,-129,-130,-129,-126,-122,-116,-109,-100,-90,-80,-69,-57,-45,-32,
	-20,-8,3,15,25,33,40,45,48,48,47,44,40,36,30,25,20,15,11,8,6,4,4
	);

	constant LUT_FIR_LPF_1k6Hz : t_lut_fir :=(
	0,1,2,3,5,7,10,13,15,17,17,16,12,7,-1,-10,-19,-29,-38,-45,-50,
	-52,-52,-49,-43,-36,-25,-14,-1,13,26,39,50,59,66,69,69,66,59,
	49,36,20,3,-14,-32,-49,-64,-77,-86,-91,-92,-88,-79,-67,-50,-30,
	-8,16,39,62,83,100,113,121,123,119,108,92,70,44,15,-17,-49,-81,
	-109,-134,-153,-165,-169,-165,-153,-132,-103,-67,-27,18,64,109,
	152,189,219,240,250,247,232,204,163,111,50,-19,-92,-166,-238,
	-304,-361,-404,-430,-437,-422,-383,-319,-230,-117,19,175,348,
	534,729,927,1123,1313,1490,1649,1787,1898,1980,2030,2047,2030,
	1980,1898,1787,1649,1490,1313,1123,927,729,534,348,175,19,-117,
	-230,-319,-383,-422,-437,-430,-404,-361,-304,-238,-166,-92,-19,
	50,111,163,204,232,247,250,240,219,189,152,109,64,18,-27,-67,-103,
	-132,-153,-165,-169,-165,-153,-134,-109,-81,-49,-17,15,44,70,92,
	108,119,123,121,113,100,83,62,39,16,-8,-30,-50,-67,-79,-88,-92,
	-91,-86,-77,-64,-49,-32,-14,3,20,36,49,59,66,69,69,66,59,50,39,
	26,13,-1,-14,-25,-36,-43,-49,-52,-52,-50,-45,-38,-29,-19,-10,-1,
	7,12,16,17,17,15,13,10,7,5,3,2,1,0
	);

	constant LUT_DELAY_MID : t_lut_fir :=(
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,32767,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	);

    constant LUT_FIR_BPF_E2 : t_lut_fir :=(
    227,258,290,324,359,396,436,478,523,571,623,679,739,803,872,945,1024,1108,1198,1294,1396,1504,1618,1740,1868,2003,2145,2295,2452,2617,2790,2970,3158,3355,3559,3772,3992,4221,4458,4703,4957,5219,5488,5766,6052,6346,6648,6957,7275,7599,7931,8271,8617,8971,9331,9697,10070,10449,10834,11224,11620,12021,12427,12837,13252,13670,14092,14518,14946,15378,15811,16247,16684,17122,17561,18001,18441,18881,19321,19759,20196,20632,21065,21496,21924,22348,22769,23186,23599,24007,24410,24807,25198,25583,25961,26333,26696,27053,27401,27741,28072,28394,28706,29009,29302,29585,29857,30119,30369,30608,30836,31052,31256,31447,31626,31793,31947,32088,32217,32332,32433,32522,32597,32658,32706,32740,32761,32768,32761,32740,32706,32658,32597,32522,32433,32332,32217,32088,31947,31793,31626,31447,31256,31052,30836,30608,30369,30119,29857,29585,29302,29009,28706,28394,28072,27741,27401,27053,26696,26333,25961,25583,25198,24807,24410,24007,23599,23186,22769,22348,21924,21496,21065,20632,20196,19759,19321,18881,18441,18001,17561,17122,16684,16247,15811,15378,14946,14518,14092,13670,13252,12837,12427,12021,11620,11224,10834,10449,10070,9697,9331,8971,8617,8271,7931,7599,7275,6957,6648,6346,6052,5766,5488,5219,4957,4703,4458,4221,3992,3772,3559,3355,3158,2970,2790,2617,2452,2295,2145,2003,1868,1740,1618,1504,1396,1294,1198,1108,1024,945,872,803,739,679,623,571,523,478,436,396,359,324,290,258,227
	);

	constant LUT_FIR_BPF_A2 : t_lut_fir :=(
    -1067,-1032,-999,-969,-941,-915,-891,-868,-845,-823,-800,-777,-752,-726,-699,-669,-636,-600,-560,-517,-469,-416,-358,-295,-225,-150,-68,20,117,221,332,452,581,718,864,1019,1183,1357,1541,1734,1938,2151,2375,2609,2854,3109,3374,3650,3937,4233,4540,4858,5185,5523,5870,6228,6595,6971,7357,7751,8155,8566,8986,9414,9850,10293,10743,11199,11662,12130,12604,13082,13565,14053,14544,15038,15534,16033,16534,17036,17539,18042,18544,19046,19546,20044,20540,21033,21522,22007,22488,22963,23433,23897,24353,24803,25245,25678,26103,26518,26924,27319,27704,28078,28440,28790,29127,29452,29763,30061,30344,30614,30869,31108,31333,31542,31735,31913,32074,32218,32346,32458,32552,32630,32690,32733,32759,32768,32759,32733,32690,32630,32552,32458,32346,32218,32074,31913,31735,31542,31333,31108,30869,30614,30344,30061,29763,29452,29127,28790,28440,28078,27704,27319,26924,26518,26103,25678,25245,24803,24353,23897,23433,22963,22488,22007,21522,21033,20540,20044,19546,19046,18544,18042,17539,17036,16534,16033,15534,15038,14544,14053,13565,13082,12604,12130,11662,11199,10743,10293,9850,9414,8986,8566,8155,7751,7357,6971,6595,6228,5870,5523,5185,4858,4540,4233,3937,3650,3374,3109,2854,2609,2375,2151,1938,1734,1541,1357,1183,1019,864,718,581,452,332,221,117,20,-68,-150,-225,-295,-358,-416,-469,-517,-560,-600,-636,-669,-699,-726,-752,-777,-800,-823,-845,-868,-891,-915,-941,-969,-999,-1032,-1067
	);

	constant LUT_FIR_BPF_D3 : t_lut_fir :=(
    -2300,-2278,-2262,-2252,-2249,-2252,-2260,-2274,-2292,-2314,-2340,-2369,-2401,-2436,-2472,-2509,-2548,-2586,-2624,-2661,-2697,-2731,-2762,-2790,-2814,-2833,-2848,-2857,-2860,-2856,-2846,-2827,-2800,-2765,-2720,-2665,-2600,-2524,-2437,-2339,-2228,-2105,-1970,-1821,-1659,-1484,-1294,-1091,-873,-641,-394,-132,143,435,741,1062,1398,1748,2114,2493,2887,3295,3717,4153,4602,5063,5538,6024,6523,7033,7553,8084,8625,9175,9734,10301,10875,11456,12044,12637,13234,13836,14441,15048,15657,16267,16878,17488,18096,18702,19306,19905,20500,21089,21672,22248,22816,23375,23925,24464,24992,25509,26013,26504,26980,27442,27889,28319,28733,29129,29508,29868,30209,30531,30832,31113,31373,31612,31829,32025,32198,32348,32476,32581,32662,32721,32756,32768,32756,32721,32662,32581,32476,32348,32198,32025,31829,31612,31373,31113,30832,30531,30209,29868,29508,29129,28733,28319,27889,27442,26980,26504,26013,25509,24992,24464,23925,23375,22816,22248,21672,21089,20500,19905,19306,18702,18096,17488,16878,16267,15657,15048,14441,13836,13234,12637,12044,11456,10875,10301,9734,9175,8625,8084,7553,7033,6523,6024,5538,5063,4602,4153,3717,3295,2887,2493,2114,1748,1398,1062,741,435,143,-132,-394,-641,-873,-1091,-1294,-1484,-1659,-1821,-1970,-2105,-2228,-2339,-2437,-2524,-2600,-2665,-2720,-2765,-2800,-2827,-2846,-2856,-2860,-2857,-2848,-2833,-2814,-2790,-2762,-2731,-2697,-2661,-2624,-2586,-2548,-2509,-2472,-2436,-2401,-2369,-2340,-2314,-2292,-2274,-2260,-2252,-2249,-2252,-2262,-2278,-2300
	);

	constant LUT_FIR_BPF_G3 : t_lut_fir :=(
    -2409,-2441,-2480,-2526,-2580,-2640,-2708,-2784,-2867,-2958,-3055,-3160,-3272,-3391,-3515,-3646,-3783,-3924,-4071,-4222,-4376,-4534,-4693,-4855,-5018,-5181,-5344,-5506,-5666,-5823,-5977,-6126,-6270,-6408,-6539,-6662,-6776,-6881,-6975,-7058,-7128,-7186,-7229,-7258,-7271,-7268,-7248,-7210,-7154,-7078,-6983,-6868,-6732,-6574,-6395,-6194,-5970,-5724,-5455,-5162,-4846,-4507,-4145,-3759,-3350,-2918,-2463,-1985,-1485,-964,-421,142,727,1331,1954,2595,3254,3930,4621,5328,6048,6781,7525,8281,9046,9819,10599,11385,12175,12969,13765,14561,15356,16150,16939,17724,18503,19273,20035,20786,21525,22251,22963,23658,24336,24996,25636,26256,26853,27426,27976,28500,28997,29468,29910,30322,30705,31057,31378,31666,31922,32145,32335,32490,32611,32698,32750,32768,32750,32698,32611,32490,32335,32145,31922,31666,31378,31057,30705,30322,29910,29468,28997,28500,27976,27426,26853,26256,25636,24996,24336,23658,22963,22251,21525,20786,20035,19273,18503,17724,16939,16150,15356,14561,13765,12969,12175,11385,10599,9819,9046,8281,7525,6781,6048,5328,4621,3930,3254,2595,1954,1331,727,142,-421,-964,-1485,-1985,-2463,-2918,-3350,-3759,-4145,-4507,-4846,-5162,-5455,-5724,-5970,-6194,-6395,-6574,-6732,-6868,-6983,-7078,-7154,-7210,-7248,-7268,-7271,-7258,-7229,-7186,-7128,-7058,-6975,-6881,-6776,-6662,-6539,-6408,-6270,-6126,-5977,-5823,-5666,-5506,-5344,-5181,-5018,-4855,-4693,-4534,-4376,-4222,-4071,-3924,-3783,-3646,-3515,-3391,-3272,-3160,-3055,-2958,-2867,-2784,-2708,-2640,-2580,-2526,-2480,-2441,-2409
	);

	constant LUT_FIR_BPF_B3 : t_lut_fir :=(
    -630,-721,-813,-909,-1009,-1113,-1222,-1338,-1460,-1589,-1726,-1871,-2025,-2187,-2359,-2541,-2732,-2933,-3143,-3364,-3594,-3833,-4082,-4339,-4605,-4878,-5159,-5447,-5740,-6039,-6342,-6649,-6958,-7268,-7579,-7889,-8198,-8503,-8804,-9099,-9387,-9667,-9937,-10196,-10442,-10675,-10892,-11093,-11276,-11440,-11582,-11703,-11801,-11874,-11922,-11942,-11935,-11899,-11833,-11737,-11609,-11448,-11255,-11028,-10768,-10473,-10143,-9778,-9379,-8945,-8475,-7972,-7433,-6861,-6256,-5618,-4948,-4247,-3516,-2756,-1967,-1152,-312,552,1439,2346,3273,4218,5178,6151,7137,8132,9134,10143,11154,12167,13179,14188,15191,16187,17172,18145,19104,20046,20969,21871,22749,23603,24429,25226,25991,26723,27421,28082,28705,29287,29829,30329,30784,31195,31560,31878,32148,32370,32544,32668,32743,32768,32743,32668,32544,32370,32148,31878,31560,31195,30784,30329,29829,29287,28705,28082,27421,26723,25991,25226,24429,23603,22749,21871,20969,20046,19104,18145,17172,16187,15191,14188,13179,12167,11154,10143,9134,8132,7137,6151,5178,4218,3273,2346,1439,552,-312,-1152,-1967,-2756,-3516,-4247,-4948,-5618,-6256,-6861,-7433,-7972,-8475,-8945,-9379,-9778,-10143,-10473,-10768,-11028,-11255,-11448,-11609,-11737,-11833,-11899,-11935,-11942,-11922,-11874,-11801,-11703,-11582,-11440,-11276,-11093,-10892,-10675,-10442,-10196,-9937,-9667,-9387,-9099,-8804,-8503,-8198,-7889,-7579,-7268,-6958,-6649,-6342,-6039,-5740,-5447,-5159,-4878,-4605,-4339,-4082,-3833,-3594,-3364,-3143,-2933,-2732,-2541,-2359,-2187,-2025,-1871,-1726,-1589,-1460,-1338,-1222,-1113,-1009,-909,-813,-721,-630
	);

	constant LUT_FIR_BPF_E4 : t_lut_fir :=(
    2494,2458,2425,2394,2364,2337,2309,2281,2251,2220,2184,2145,2099,2047,1986,1917,1836,1744,1639,1520,1386,1235,1067,881,676,450,204,-62,-351,-662,-995,-1350,-1727,-2127,-2548,-2990,-3452,-3934,-4434,-4952,-5486,-6034,-6596,-7169,-7751,-8340,-8935,-9533,-10131,-10728,-11320,-11904,-12480,-13042,-13589,-14118,-14626,-15110,-15567,-15995,-16390,-16750,-17072,-17354,-17593,-17787,-17933,-18030,-18075,-18066,-18003,-17883,-17705,-17468,-17172,-16815,-16398,-15919,-15380,-14780,-14121,-13402,-12625,-11791,-10901,-9958,-8964,-7920,-6829,-5693,-4517,-3302,-2052,-770,538,1872,3226,4597,5979,7370,8764,10157,11545,12923,14287,15633,16956,18251,19515,20743,21930,23074,24169,25213,26202,27132,28000,28803,29538,30203,30795,31313,31754,32117,32401,32604,32727,32768,32727,32604,32401,32117,31754,31313,30795,30203,29538,28803,28000,27132,26202,25213,24169,23074,21930,20743,19515,18251,16956,15633,14287,12923,11545,10157,8764,7370,5979,4597,3226,1872,538,-770,-2052,-3302,-4517,-5693,-6829,-7920,-8964,-9958,-10901,-11791,-12625,-13402,-14121,-14780,-15380,-15919,-16398,-16815,-17172,-17468,-17705,-17883,-18003,-18066,-18075,-18030,-17933,-17787,-17593,-17354,-17072,-16750,-16390,-15995,-15567,-15110,-14626,-14118,-13589,-13042,-12480,-11904,-11320,-10728,-10131,-9533,-8935,-8340,-7751,-7169,-6596,-6034,-5486,-4952,-4434,-3934,-3452,-2990,-2548,-2127,-1727,-1350,-995,-662,-351,-62,204,450,676,881,1067,1235,1386,1520,1639,1744,1836,1917,1986,2047,2099,2145,2184,2220,2251,2281,2309,2337,2364,2394,2425,2458,2494
	);
    
 	
	-------------------------------------------------------------------------------		
end package;
