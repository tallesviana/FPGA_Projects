-------------------------------------------
--    Title   
--    Description   
-- 
--

LIBRARY ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--||||||   ENTITY   ||||||--

ENTITY xxxxx IS
    GENERIC(

    );
    PORT(
        
    );
END xxxxx;

--||||||   ARCHITECTURE  ||||||--

ARCHITECTURE rtl OF xxxxx IS

BEGIN

    -->> Combination Logic

    -->> Sequential Logic

    -->> Concurrent Assignments

END rtl;