-------------------------------------------------------------------------------
-- Project     : Audio_Synth
-- Description : Constants and LUT for audio filters
--
--
-------------------------------------------------------------------------------
--
-- Change History
-- Date     |Name      |Modification
------------|----------|-------------------------------------------------------
-- 26.03.18 | dqtm     | file created for EA-999 demo
-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
-- Package  Declaration
-------------------------------------------------------------------------------
-- Include in Design of filter blocks, using  :
--   use work.audio_filter_pkg.all;
-------------------------------------------------------------------------------
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

package audio_filter_pkg is

    --constant N_CUM:					natural :=19; 			-- number of bits in phase cumulator phicum_reg
	--constant N_AUDIO :				natural := 16;			-- Audio Paralell Bus width

    -------------------------------------------------------------------------------
	-- CONSTANT & TYPES FOR FIR 
	-------------------------------------------------------------------------------
    constant N_RESOL_TAP:			natural := 32;  		-- resolution of each position on tap-line (storing MAC outputs)
    constant N_LUT:					natural := 255;  		-- length of LUT = 255
	constant N_addr_LUT:			natural := 8; 			-- number of bits to address LUT (for index)
	
    constant N_RESOL_COEFF:			natural := 16;			-- Attention: 1 bit reserved for sign, FIR-coeffs use 12-bits
															-- range : [-2^15; +(2^15)-1] = [-32768 ; +32767]
															-- but from Matlab file expect scaling fitting in the
															-- range : [-2^11; +(2^11)-1] = [-2048 ; +2047]
    subtype  t_fir_range is integer range -(2**(N_RESOL_COEFF-1)) to (2**(N_RESOL_COEFF-1))-1;
	type     t_lut_fir is array (0 to N_LUT-1) of t_fir_range;


	constant LUT_FIR_LPF_200Hz : t_lut_fir :=(
	-14,-15,-19,-25,-34,-45,-58,-73,-90,-109,-129,-149,-170,-189,-208,
	-226,-241,-253,-263,-269,-272,-273,-273,-273,-272,-270,-268,-265,-262,
	-257,-252,-247,-240,-233,-225,-216,-207,-197,-186,-174,-161,-147,-133,
	-118,-102,-85,-67,-49,-29,-9,12,33,56,79,103,128,154,180,207,235,264,
	293,322,353,384,415,447,480,513,547,580,615,649,685,720,755,791,827,
	863,900,936,972,1009,1045,1081,1118,1154,1189,1225,1260,1295,1330,
	1364,1398,1431,1464,1496,1528,1559,1589,1619,1648,1676,1703,1730,1755,
	1780,1804,1827,1848,1869,1889,1908,1925,1942,1957,1971,1984,1996,2007,
	2016,2024,2031,2037,2041,2044,2046,2047,2046,2044,2041,2037,2031,2024,
	2016,2007,1996,1984,1971,1957,1942,1925,1908,1889,1869,1848,1827,1804,
	1780,1755,1730,1703,1676,1648,1619,1589,1559,1528,1496,1464,1431,1398,
	1364,1330,1295,1260,1225,1189,1154,1118,1081,1045,1009,972,936,900,
	863,827,791,755,720,685,649,615,580,547,513,480,447,415,384,353,322,
	293,264,235,207,180,154,128,103,79,56,33,12,-9,-29,-49,-67,-85,-102,
	-118,-133,-147,-161,-174,-186,-197,-207,-216,-225,-233,-240,-247,-252,
	-257,-262,-265,-268,-270,-272,-273,-273,-273,-272,-269,-263,-253,-241,
	-226,-208,-189,-170,-149,-129,-109,-90,-73,-58,-45,-34,-25,-19,-15,-14
	);
	
	constant LUT_FIR_LPF_400Hz : t_lut_fir :=(
	8,9,11,15,21,27,35,45,55,66,77,89,99,109,118,124,129,132,132,130,125,
	119,112,104,95,86,75,64,52,40,26,12,-2,-17,-33,-49,-65,-82,-99,-116,
	-134,-151,-168,-185,-202,-219,-235,-251,-266,-281,-295,-308,-320,-330,
	-340,-349,-356,-362,-366,-369,-370,-370,-367,-363,-357,-349,-339,-327,
	-312,-296,-278,-257,-234,-209,-182,-153,-121,-88,-52,-15,25,66,110,
	155,201,250,300,351,404,458,513,569,625,683,741,799,858,917,976,1034,
	1093,1151,1208,1264,1320,1374,1428,1480,1530,1579,1626,1671,1714,1755,
	1793,1830,1863,1894,1923,1948,1971,1991,2008,2022,2033,2041,2045,2047,
	2045,2041,2033,2022,2008,1991,1971,1948,1923,1894,1863,1830,1793,1755,
	1714,1671,1626,1579,1530,1480,1428,1374,1320,1264,1208,1151,1093,1034,
	976,917,858,799,741,683,625,569,513,458,404,351,300,250,201,155,110,
	66,25,-15,-52,-88,-121,-153,-182,-209,-234,-257,-278,-296,-312,-327,
	-339,-349,-357,-363,-367,-370,-370,-369,-366,-362,-356,-349,-340,-330,
	-320,-308,-295,-281,-266,-251,-235,-219,-202,-185,-168,-151,-134,-116,
	-99,-82,-65,-49,-33,-17,-2,12,26,40,52,64,75,86,95,104,112,119,125,
	130,132,132,129,124,118,109,99,89,77,66,55,45,35,27,21,15,11,9,8
	);

	constant LUT_FIR_LPF_800Hz : t_lut_fir :=(
	4,4,6,8,11,15,20,25,30,36,40,44,47,48,48,45,40,33,25,15,3,-8,-20,
	-32,-45,-57,-69,-80,-90,-100,-109,-116,-122,-126,-129,-130,-129,
	-126,-121,-115,-106,-96,-83,-69,-54,-37,-19,0,20,41,61,82,102,122,
	140,158,174,188,199,209,216,220,220,218,213,204,192,177,158,136,
	111,84,54,22,-12,-47,-84,-121,-158,-194,-230,-264,-296,-326,-352,
	-375,-394,-408,-416,-420,-417,-408,-393,-371,-342,-306,-263,-213,
	-157,-94,-24,52,133,219,310,405,504,605,708,813,918,1023,1126,1228,
	1327,1422,1513,1599,1679,1753,1819,1878,1929,1971,2004,2028,2042,
	2047,2042,2028,2004,1971,1929,1878,1819,1753,1679,1599,1513,1422,
	1327,1228,1126,1023,918,813,708,605,504,405,310,219,133,52,-24,-94,
	-157,-213,-263,-306,-342,-371,-393,-408,-417,-420,-416,-408,-394,
	-375,-352,-326,-296,-264,-230,-194,-158,-121,-84,-47,-12,22,54,84,
	111,136,158,177,192,204,213,218,220,220,216,209,199,188,174,158,
	140,122,102,82,61,41,20,0,-19,-37,-54,-69,-83,-96,-106,-115,-121,
	-126,-129,-130,-129,-126,-122,-116,-109,-100,-90,-80,-69,-57,-45,-32,
	-20,-8,3,15,25,33,40,45,48,48,47,44,40,36,30,25,20,15,11,8,6,4,4
	);

	constant LUT_FIR_LPF_1k6Hz : t_lut_fir :=(
	0,1,2,3,5,7,10,13,15,17,17,16,12,7,-1,-10,-19,-29,-38,-45,-50,
	-52,-52,-49,-43,-36,-25,-14,-1,13,26,39,50,59,66,69,69,66,59,
	49,36,20,3,-14,-32,-49,-64,-77,-86,-91,-92,-88,-79,-67,-50,-30,
	-8,16,39,62,83,100,113,121,123,119,108,92,70,44,15,-17,-49,-81,
	-109,-134,-153,-165,-169,-165,-153,-132,-103,-67,-27,18,64,109,
	152,189,219,240,250,247,232,204,163,111,50,-19,-92,-166,-238,
	-304,-361,-404,-430,-437,-422,-383,-319,-230,-117,19,175,348,
	534,729,927,1123,1313,1490,1649,1787,1898,1980,2030,2047,2030,
	1980,1898,1787,1649,1490,1313,1123,927,729,534,348,175,19,-117,
	-230,-319,-383,-422,-437,-430,-404,-361,-304,-238,-166,-92,-19,
	50,111,163,204,232,247,250,240,219,189,152,109,64,18,-27,-67,-103,
	-132,-153,-165,-169,-165,-153,-134,-109,-81,-49,-17,15,44,70,92,
	108,119,123,121,113,100,83,62,39,16,-8,-30,-50,-67,-79,-88,-92,
	-91,-86,-77,-64,-49,-32,-14,3,20,36,49,59,66,69,69,66,59,50,39,
	26,13,-1,-14,-25,-36,-43,-49,-52,-52,-50,-45,-38,-29,-19,-10,-1,
	7,12,16,17,17,15,13,10,7,5,3,2,1,0
	);

	constant LUT_DELAY_MID : t_lut_fir :=(
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,32767,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	);

	constant LUT_FIR_BPF_E2_v2 : t_lut_fir :=(
	227,258,290,324,359,396,436,478,523,571,623,679,739,803,871,945,1024,1108,1198,1294,1396,1504,1618,1740,1868,2003,2145,2295,2452,2617,2790,2970,3158,3355,3559,3771,3992,4221,4458,4703,4957,5218,5488,5766,6052,6346,6648,6957,7274,7599,7931,8271,8617,8970,9330,9697,10070,10449,10834,11224,11620,12021,12427,12837,13251,13670,14092,14517,14946,15377,15811,16246,16683,17122,17561,18001,18441,18881,19320,19759,20196,20631,21064,21495,21923,22348,22769,23186,23598,24006,24409,24806,25197,25582,25960,26332,26696,27052,27400,27740,28071,28393,28705,29008,29301,29584,29856,30118,30368,30607,30835,31051,31255,31446,31626,31792,31946,32087,32216,32331,32432,32521,32596,32657,32705,32739,32760,32767,32760,32739,32705,32657,32596,32521,32432,32331,32216,32087,31946,31792,31626,31446,31255,31051,30835,30607,30368,30118,29856,29584,29301,29008,28705,28393,28071,27740,27400,27052,26696,26332,25960,25582,25197,24806,24409,24006,23598,23186,22769,22348,21923,21495,21064,20631,20196,19759,19320,18881,18441,18001,17561,17122,16683,16246,15811,15377,14946,14517,14092,13670,13251,12837,12427,12021,11620,11224,10834,10449,10070,9697,9330,8970,8617,8271,7931,7599,7274,6957,6648,6346,6052,5766,5488,5218,4957,4703,4458,4221,3992,3771,3559,3355,3158,2970,2790,2617,2452,2295,2145,2003,1868,1740,1618,1504,1396,1294,1198,1108,1024,945,871,803,739,679,623,571,523,478,436,396,359,324,290,258,227
	);

	constant LUT_FIR_BPF_E4_v2 : t_lut_fir :=(
	2494,2458,2425,2394,2364,2336,2309,2281,2251,2220,2184,2145,2099,2047,1986,1917,1836,1744,1639,1520,1386,1235,1067,881,676,450,204,-62,-351,-662,-995,-1350,-1727,-2127,-2548,-2990,-3452,-3934,-4434,-4952,-5486,-6034,-6596,-7168,-7751,-8340,-8935,-9533,-10131,-10727,-11319,-11904,-12479,-13042,-13589,-14118,-14626,-15110,-15567,-15994,-16389,-16749,-17072,-17354,-17593,-17786,-17932,-18029,-18074,-18066,-18002,-17882,-17704,-17468,-17171,-16814,-16397,-15919,-15380,-14780,-14120,-13401,-12624,-11790,-10901,-9958,-8963,-7919,-6828,-5693,-4517,-3302,-2052,-770,538,1872,3226,4597,5979,7369,8763,10157,11545,12923,14287,15633,16955,18251,19514,20742,21930,23073,24169,25213,26201,27131,27999,28802,29537,30202,30794,31312,31753,32116,32400,32603,32726,32767,32726,32603,32400,32116,31753,31312,30794,30202,29537,28802,27999,27131,26201,25213,24169,23073,21930,20742,19514,18251,16955,15633,14287,12923,11545,10157,8763,7369,5979,4597,3226,1872,538,-770,-2052,-3302,-4517,-5693,-6828,-7919,-8963,-9958,-10901,-11790,-12624,-13401,-14120,-14780,-15380,-15919,-16397,-16814,-17171,-17468,-17704,-17882,-18002,-18066,-18074,-18029,-17932,-17786,-17593,-17354,-17072,-16749,-16389,-15994,-15567,-15110,-14626,-14118,-13589,-13042,-12479,-11904,-11319,-10727,-10131,-9533,-8935,-8340,-7751,-7168,-6596,-6034,-5486,-4952,-4434,-3934,-3452,-2990,-2548,-2127,-1727,-1350,-995,-662,-351,-62,204,450,676,881,1067,1235,1386,1520,1639,1744,1836,1917,1986,2047,2099,2145,2184,2220,2251,2281,2309,2336,2364,2394,2425,2458,2494
	);

	constant LUT_FIR_LPF_100Hz_v2 : t_lut_fir :=(
	1407,1426,1449,1478,1512,1552,1597,1649,1706,1769,1839,1915,1997,2086,2182,2284,2394,2510,2633,2764,2901,3046,3198,3358,3524,3699,3880,4069,4265,4469,4680,4898,5123,5356,5596,5843,6098,6359,6627,6902,7184,7472,7767,8068,8376,8690,9009,9335,9666,10003,10345,10692,11044,11400,11762,12127,12497,12870,13248,13628,14012,14399,14788,15180,15574,15970,16367,16766,17166,17567,17968,18370,18771,19172,19573,19973,20371,20768,21163,21556,21946,22334,22719,23100,23478,23852,24222,24587,24948,25304,25654,25999,26337,26670,26996,27316,27628,27934,28232,28522,28805,29079,29345,29602,29851,30091,30321,30542,30753,30955,31147,31328,31500,31661,31811,31951,32080,32198,32306,32402,32487,32561,32624,32675,32715,32744,32761,32767,32761,32744,32715,32675,32624,32561,32487,32402,32306,32198,32080,31951,31811,31661,31500,31328,31147,30955,30753,30542,30321,30091,29851,29602,29345,29079,28805,28522,28232,27934,27628,27316,26996,26670,26337,25999,25654,25304,24948,24587,24222,23852,23478,23100,22719,22334,21946,21556,21163,20768,20371,19973,19573,19172,18771,18370,17968,17567,17166,16766,16367,15970,15574,15180,14788,14399,14012,13628,13248,12870,12497,12127,11762,11400,11044,10692,10345,10003,9666,9335,9009,8690,8376,8068,7767,7472,7184,6902,6627,6359,6098,5843,5596,5356,5123,4898,4680,4469,4265,4069,3880,3699,3524,3358,3198,3046,2901,2764,2633,2510,2394,2284,2182,2086,1997,1915,1839,1769,1706,1649,1597,1552,1512,1478,1449,1426,1407
	);

	constant LUT_FIR_LPF_200Hz_v2 : t_lut_fir :=(
	-332,-317,-302,-287,-273,-258,-243,-228,-212,-195,-176,-156,-135,-111,-85,-56,-25,8,46,88,134,184,239,298,363,433,509,592,680,776,878,987,1104,1229,1361,1502,1651,1809,1976,2151,2336,2530,2734,2947,3171,3404,3647,3900,4163,4436,4719,5012,5316,5629,5953,6286,6630,6983,7345,7717,8098,8488,8887,9294,9710,10134,10565,11004,11450,11903,12361,12826,13297,13772,14253,14737,15225,15717,16211,16708,17207,17706,18207,18708,19208,19707,20205,20701,21195,21685,22171,22653,23130,23601,24067,24526,24977,25421,25856,26283,26700,27107,27503,27889,28263,28624,28974,29310,29633,29943,30237,30518,30783,31033,31267,31485,31687,31872,32041,32192,32326,32442,32541,32622,32685,32730,32757,32767,32757,32730,32685,32622,32541,32442,32326,32192,32041,31872,31687,31485,31267,31033,30783,30518,30237,29943,29633,29310,28974,28624,28263,27889,27503,27107,26700,26283,25856,25421,24977,24526,24067,23601,23130,22653,22171,21685,21195,20701,20205,19707,19208,18708,18207,17706,17207,16708,16211,15717,15225,14737,14253,13772,13297,12826,12361,11903,11450,11004,10565,10134,9710,9294,8887,8488,8098,7717,7345,6983,6630,6286,5953,5629,5316,5012,4719,4436,4163,3900,3647,3404,3171,2947,2734,2530,2336,2151,1976,1809,1651,1502,1361,1229,1104,987,878,776,680,592,509,433,363,298,239,184,134,88,46,8,-25,-56,-85,-111,-135,-156,-176,-195,-212,-228,-243,-258,-273,-287,-302,-317,-332
	);

	constant LUT_FIR_LPF_400Hz_v2 : t_lut_fir :=(
	295,285,276,265,255,244,232,219,205,190,173,154,133,110,85,56,25,-8,-46,-88,-133,-183,-236,-293,-355,-421,-492,-567,-646,-729,-816,-907,-1001,-1099,-1200,-1303,-1409,-1516,-1624,-1733,-1842,-1950,-2056,-2160,-2262,-2359,-2451,-2538,-2618,-2691,-2754,-2809,-2852,-2884,-2902,-2907,-2897,-2872,-2829,-2768,-2688,-2588,-2467,-2325,-2160,-1972,-1760,-1523,-1261,-974,-660,-319,47,441,862,1310,1785,2287,2815,3369,3948,4552,5180,5831,6505,7200,7914,8648,9399,10166,10948,11743,12549,13364,14188,15017,15849,16684,17519,18351,19180,20001,20814,21617,22407,23181,23939,24678,25395,26089,26758,27400,28014,28596,29146,29662,30143,30587,30993,31359,31685,31969,32211,32410,32566,32677,32744,32767,32744,32677,32566,32410,32211,31969,31685,31359,30993,30587,30143,29662,29146,28596,28014,27400,26758,26089,25395,24678,23939,23181,22407,21617,20814,20001,19180,18351,17519,16684,15849,15017,14188,13364,12549,11743,10948,10166,9399,8648,7914,7200,6505,5831,5180,4552,3948,3369,2815,2287,1785,1310,862,441,47,-319,-660,-974,-1261,-1523,-1760,-1972,-2160,-2325,-2467,-2588,-2688,-2768,-2829,-2872,-2897,-2907,-2902,-2884,-2852,-2809,-2754,-2691,-2618,-2538,-2451,-2359,-2262,-2160,-2056,-1950,-1842,-1733,-1624,-1516,-1409,-1303,-1200,-1099,-1001,-907,-816,-729,-646,-567,-492,-421,-355,-293,-236,-183,-133,-88,-46,-8,25,56,85,110,133,154,173,190,205,219,232,244,255,265,276,285,295
	);
	-------------------------------------------------------------------------------		
end package;
