-------------------------------------------------------------------------------
-- Project     : Audio_Synth
-- Description : Constants and LUT for audio filters
--
--
-------------------------------------------------------------------------------
--
-- Change History
-- Date     |Name      |Modification
------------|----------|-------------------------------------------------------
-- 26.03.18 | dqtm     | file created for EA-999 demo
-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
-- Package  Declaration
-------------------------------------------------------------------------------
-- Include in Design of filter blocks, using  :
--   use work.audio_filter_pkg.all;
-------------------------------------------------------------------------------
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

package audio_filter_pkg is

    --constant N_CUM:					natural :=19; 			-- number of bits in phase cumulator phicum_reg
	--constant N_AUDIO :				natural := 16;			-- Audio Paralell Bus width

    -------------------------------------------------------------------------------
	-- CONSTANT & TYPES FOR FIR 
	-------------------------------------------------------------------------------
    constant N_RESOL_TAP:			natural := 32;  		-- resolution of each position on tap-line (storing MAC outputs)
    constant N_LUT:					natural := 255;  		-- length of LUT = 255
	constant N_addr_LUT:			natural := 8; 			-- number of bits to address LUT (for index)
	
    constant N_RESOL_COEFF:			natural := 16;			-- Attention: 1 bit reserved for sign, FIR-coeffs use 12-bits
															-- range : [-2^15; +(2^15)-1] = [-32768 ; +32767]
															-- but from Matlab file expect scaling fitting in the
															-- range : [-2^11; +(2^11)-1] = [-2048 ; +2047]
    subtype  t_fir_range is integer range -(2**(N_RESOL_COEFF-1)) to (2**(N_RESOL_COEFF-1))-1;
	type     t_lut_fir is array (0 to N_LUT-1) of t_fir_range;


	constant LUT_FIR_LPF_200Hz : t_lut_fir :=(
	-14,-15,-19,-25,-34,-45,-58,-73,-90,-109,-129,-149,-170,-189,-208,
	-226,-241,-253,-263,-269,-272,-273,-273,-273,-272,-270,-268,-265,-262,
	-257,-252,-247,-240,-233,-225,-216,-207,-197,-186,-174,-161,-147,-133,
	-118,-102,-85,-67,-49,-29,-9,12,33,56,79,103,128,154,180,207,235,264,
	293,322,353,384,415,447,480,513,547,580,615,649,685,720,755,791,827,
	863,900,936,972,1009,1045,1081,1118,1154,1189,1225,1260,1295,1330,
	1364,1398,1431,1464,1496,1528,1559,1589,1619,1648,1676,1703,1730,1755,
	1780,1804,1827,1848,1869,1889,1908,1925,1942,1957,1971,1984,1996,2007,
	2016,2024,2031,2037,2041,2044,2046,2047,2046,2044,2041,2037,2031,2024,
	2016,2007,1996,1984,1971,1957,1942,1925,1908,1889,1869,1848,1827,1804,
	1780,1755,1730,1703,1676,1648,1619,1589,1559,1528,1496,1464,1431,1398,
	1364,1330,1295,1260,1225,1189,1154,1118,1081,1045,1009,972,936,900,
	863,827,791,755,720,685,649,615,580,547,513,480,447,415,384,353,322,
	293,264,235,207,180,154,128,103,79,56,33,12,-9,-29,-49,-67,-85,-102,
	-118,-133,-147,-161,-174,-186,-197,-207,-216,-225,-233,-240,-247,-252,
	-257,-262,-265,-268,-270,-272,-273,-273,-273,-272,-269,-263,-253,-241,
	-226,-208,-189,-170,-149,-129,-109,-90,-73,-58,-45,-34,-25,-19,-15,-14
	);
	
	constant LUT_FIR_LPF_400Hz : t_lut_fir :=(
	8,9,11,15,21,27,35,45,55,66,77,89,99,109,118,124,129,132,132,130,125,
	119,112,104,95,86,75,64,52,40,26,12,-2,-17,-33,-49,-65,-82,-99,-116,
	-134,-151,-168,-185,-202,-219,-235,-251,-266,-281,-295,-308,-320,-330,
	-340,-349,-356,-362,-366,-369,-370,-370,-367,-363,-357,-349,-339,-327,
	-312,-296,-278,-257,-234,-209,-182,-153,-121,-88,-52,-15,25,66,110,
	155,201,250,300,351,404,458,513,569,625,683,741,799,858,917,976,1034,
	1093,1151,1208,1264,1320,1374,1428,1480,1530,1579,1626,1671,1714,1755,
	1793,1830,1863,1894,1923,1948,1971,1991,2008,2022,2033,2041,2045,2047,
	2045,2041,2033,2022,2008,1991,1971,1948,1923,1894,1863,1830,1793,1755,
	1714,1671,1626,1579,1530,1480,1428,1374,1320,1264,1208,1151,1093,1034,
	976,917,858,799,741,683,625,569,513,458,404,351,300,250,201,155,110,
	66,25,-15,-52,-88,-121,-153,-182,-209,-234,-257,-278,-296,-312,-327,
	-339,-349,-357,-363,-367,-370,-370,-369,-366,-362,-356,-349,-340,-330,
	-320,-308,-295,-281,-266,-251,-235,-219,-202,-185,-168,-151,-134,-116,
	-99,-82,-65,-49,-33,-17,-2,12,26,40,52,64,75,86,95,104,112,119,125,
	130,132,132,129,124,118,109,99,89,77,66,55,45,35,27,21,15,11,9,8
	);

	constant LUT_FIR_LPF_800Hz : t_lut_fir :=(
	4,4,6,8,11,15,20,25,30,36,40,44,47,48,48,45,40,33,25,15,3,-8,-20,
	-32,-45,-57,-69,-80,-90,-100,-109,-116,-122,-126,-129,-130,-129,
	-126,-121,-115,-106,-96,-83,-69,-54,-37,-19,0,20,41,61,82,102,122,
	140,158,174,188,199,209,216,220,220,218,213,204,192,177,158,136,
	111,84,54,22,-12,-47,-84,-121,-158,-194,-230,-264,-296,-326,-352,
	-375,-394,-408,-416,-420,-417,-408,-393,-371,-342,-306,-263,-213,
	-157,-94,-24,52,133,219,310,405,504,605,708,813,918,1023,1126,1228,
	1327,1422,1513,1599,1679,1753,1819,1878,1929,1971,2004,2028,2042,
	2047,2042,2028,2004,1971,1929,1878,1819,1753,1679,1599,1513,1422,
	1327,1228,1126,1023,918,813,708,605,504,405,310,219,133,52,-24,-94,
	-157,-213,-263,-306,-342,-371,-393,-408,-417,-420,-416,-408,-394,
	-375,-352,-326,-296,-264,-230,-194,-158,-121,-84,-47,-12,22,54,84,
	111,136,158,177,192,204,213,218,220,220,216,209,199,188,174,158,
	140,122,102,82,61,41,20,0,-19,-37,-54,-69,-83,-96,-106,-115,-121,
	-126,-129,-130,-129,-126,-122,-116,-109,-100,-90,-80,-69,-57,-45,-32,
	-20,-8,3,15,25,33,40,45,48,48,47,44,40,36,30,25,20,15,11,8,6,4,4
	);

	constant LUT_FIR_LPF_1k6Hz : t_lut_fir :=(
	0,1,2,3,5,7,10,13,15,17,17,16,12,7,-1,-10,-19,-29,-38,-45,-50,
	-52,-52,-49,-43,-36,-25,-14,-1,13,26,39,50,59,66,69,69,66,59,
	49,36,20,3,-14,-32,-49,-64,-77,-86,-91,-92,-88,-79,-67,-50,-30,
	-8,16,39,62,83,100,113,121,123,119,108,92,70,44,15,-17,-49,-81,
	-109,-134,-153,-165,-169,-165,-153,-132,-103,-67,-27,18,64,109,
	152,189,219,240,250,247,232,204,163,111,50,-19,-92,-166,-238,
	-304,-361,-404,-430,-437,-422,-383,-319,-230,-117,19,175,348,
	534,729,927,1123,1313,1490,1649,1787,1898,1980,2030,2047,2030,
	1980,1898,1787,1649,1490,1313,1123,927,729,534,348,175,19,-117,
	-230,-319,-383,-422,-437,-430,-404,-361,-304,-238,-166,-92,-19,
	50,111,163,204,232,247,250,240,219,189,152,109,64,18,-27,-67,-103,
	-132,-153,-165,-169,-165,-153,-134,-109,-81,-49,-17,15,44,70,92,
	108,119,123,121,113,100,83,62,39,16,-8,-30,-50,-67,-79,-88,-92,
	-91,-86,-77,-64,-49,-32,-14,3,20,36,49,59,66,69,69,66,59,50,39,
	26,13,-1,-14,-25,-36,-43,-49,-52,-52,-50,-45,-38,-29,-19,-10,-1,
	7,12,16,17,17,15,13,10,7,5,3,2,1,0
	);

	constant LUT_DELAY_MID : t_lut_fir :=(
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,32767,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	);

 	
	-------------------------------------------------------------------------------		
end package;
